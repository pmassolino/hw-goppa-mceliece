----------------------------------------------------------------------------------
-- Company: LARC - Escola Politecnica - University of Sao Paulo
-- Engineer: Pedro Maat C. Massolino
-- 
-- Create Date:    05/12/2012 
-- Design Name:    Controller_Solving_Key_Equation_1_v2
-- Module Name:    Controller_Solving_Key_Equation_1_v2
-- Project Name:   McEliece QD-Goppa Decoder
-- Target Devices: Any
-- Tool versions:  Xilinx ISE 13.3 WebPack
--
-- Description: 
-- 
-- The 2nd step in Goppa Code Decoding.
--
-- This is a state machine circuit that controls solving_key_equation_1_v2.
-- This state machine have 3 phases: first phase variable initialization,
-- second computation of polynomial sigma, third step writing the polynomial sigma
-- on a specific memory position.
--
-- This is the second circuit version. It is a non pipeline version of the algorithm, 
-- each coefficient takes more than 1 cycle to be computed.
-- A more optimized pipelined version was made called solving_key_equation_2
--
-- Dependencies: 
--
-- VHDL-93
--
-- Revision: 
-- Revision 1.0
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity controller_solving_key_equation_1_v2 is
	Port(
		clk : in STD_LOGIC;
		rst : in STD_LOGIC;
		FB_equal_zero : in STD_LOGIC;
		i_equal_zero : in STD_LOGIC;
		i_minus_j_less_than_zero : in STD_LOGIC;
		degree_G_less_equal_final_degree : in STD_LOGIC;
		degree_F_less_than_degree_G : in STD_LOGIC;
		degree_B_equal_degree_C_plus_j : in STD_LOGIC;
		degree_B_less_than_degree_C_plus_j : in STD_LOGIC;
		reg_looking_degree_q : in STD_LOGIC_VECTOR(0 downto 0);
		key_equation_found : out STD_LOGIC;
		signal_inv : out STD_LOGIC;
		sel_new_value_inv : out STD_LOGIC;
		write_enable_FB : out STD_LOGIC;
		write_enable_GC : out STD_LOGIC;
		sel_base_mul : out STD_LOGIC;
		reg_h_ce : out STD_LOGIC;
		ctr_i_ce : out STD_LOGIC;
		ctr_i_load : out STD_LOGIC;
		ctr_i_rst : out STD_LOGIC;
		sel_ctr_i_rst_value : out STD_LOGIC;
		sel_ctr_i_d : out STD_LOGIC;
		reg_j_ce : out STD_LOGIC;
		reg_j_rst : out STD_LOGIC;
		reg_FB_ce : out STD_LOGIC;
		reg_FB_rst : out STD_LOGIC;
		sel_reg_FB : out STD_LOGIC;
		sel_load_new_value_FB : out STD_LOGIC;
		reg_GC_ce : out STD_LOGIC;
		reg_GC_rst : out STD_LOGIC;
		sel_reg_GC : out STD_LOGIC;
		ctr_degree_F_ce : out STD_LOGIC;
		ctr_degree_F_load : out STD_LOGIC;
		ctr_degree_F_rst : out STD_LOGIC;
		reg_degree_G_ce : out STD_LOGIC;
		reg_degree_G_rst : out STD_LOGIC;
		ctr_degree_B_ce : out STD_LOGIC;
		ctr_degree_B_load : out STD_LOGIC;
		ctr_degree_B_rst : out STD_LOGIC;
		sel_ctr_degree_B : out STD_LOGIC;
		reg_degree_C_ce : out STD_LOGIC;
		reg_degree_C_rst : out STD_LOGIC;
		reg_looking_degree_d : out STD_LOGIC_VECTOR(0 downto 0);
		reg_looking_degree_ce : out STD_LOGIC;
		reg_swap_ce : out STD_LOGIC;
		reg_swap_rst : out STD_LOGIC;
		sel_address_FB : out STD_LOGIC;
		sel_address_GC : out STD_LOGIC;
		ctr_address_FB_ce : out STD_LOGIC;
		ctr_address_FB_load : out STD_LOGIC;
		ctr_address_GC_ce : out STD_LOGIC;
		ctr_address_GC_load : out STD_LOGIC;
		BC_calculation : out STD_LOGIC;
		enable_external_swap : out STD_LOGIC
	);
end controller_solving_key_equation_1_v2;

architecture Behavioral of controller_solving_key_equation_1_v2 is

type State is (reset, load_counter, store_G2t, load_first_inv, send_first_inv, prepare_load_F_store_G, load_F_store_G, wait_F, prepare_store_B_C, store_B_C, last_store_B_C, swap_F_G_B_C, prepare_load_j, load_j, load_first_G_first_F, load_h, prepare_load_F_G, load_F_G, mult_add_F_G, store_F, finalize_i, prepare_i, prepare_load_B_C, load_B_C, mult_add_B_C, store_B, prepare_final_swap, preparel_swap_address, prepare_load_sigma, load_sigma, store_sigma, final); 
signal actual_state, next_state : State; 

begin

Clock: process (clk)
begin
	if (clk'event and clk = '1') then
		if (rst = '1') then
			actual_state <= reset;
		else
			actual_state <= next_state;
		end if;        
	end if;
end process;

Output: process(actual_state, FB_equal_zero, i_equal_zero, i_minus_j_less_than_zero, degree_G_less_equal_final_degree, degree_F_less_than_degree_G,	degree_B_equal_degree_C_plus_j, degree_B_less_than_degree_C_plus_j, reg_looking_degree_q)
begin
	case (actual_state) is
		when reset =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= '1';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '1';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '1';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '1';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_counter =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= '1';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '1';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '1';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '1';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '1';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= '1';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when store_G2t =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';			
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= '1';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '1';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '1';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "1";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_first_inv =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';			
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when send_first_inv =>
			key_equation_found <= '0';
			signal_inv <= '1';
			sel_new_value_inv <= '1';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';			
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_F_store_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_F_store_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when wait_F =>
			if(i_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';				
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '1';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			elsif(reg_looking_degree_q(0) = '1' and FB_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '1';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when prepare_store_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';				
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when store_B_C =>
			if(i_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '1';
				sel_base_mul <= '0';
				reg_h_ce <= '0';				
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '1';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '1';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '1';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when last_store_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '1';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '1';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			BC_calculation <= '1';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			enable_external_swap <= '1';
		when swap_F_G_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '1';
			ctr_degree_F_load <= '1';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '1';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '1';
			ctr_degree_B_load <= '1';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '1';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '1';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_j =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_rst <= '0';
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '1';
			sel_address_GC <= '1';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_j =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '1';
			ctr_i_load <= '1';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '1';
			reg_j_ce <= '1';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '1';
			sel_address_GC <= '1';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_first_G_first_F =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '1';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_h =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '1';
			reg_h_ce <= '1';	
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "1";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_F_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_F_G =>
			if(i_minus_j_less_than_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '1';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when mult_add_F_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '1';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when store_F =>
			if(i_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_load_new_value_FB <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			elsif(reg_looking_degree_q(0) = '1') then
				if(FB_equal_zero = '1') then
					key_equation_found <= '0';
					signal_inv <= '0';
					sel_new_value_inv <= '0';
					write_enable_FB <= '1';
					write_enable_GC <= '0';
					sel_base_mul <= '0';
					reg_h_ce <= '0';
					ctr_i_ce <= '1';
					ctr_i_load <= '0';
					ctr_i_rst <= '0';
					sel_ctr_i_rst_value <= '0';
					sel_ctr_i_d <= '0';
					reg_j_ce <= '0';
					reg_j_rst <= '0';
					reg_FB_ce <= '0';
					reg_FB_rst <= '0';
					sel_reg_FB <= '0';
					sel_load_new_value_FB <= '0';
					reg_GC_ce <= '0';
					reg_GC_rst <= '0';
					sel_reg_GC <= '0';
					ctr_degree_F_ce <= '1';
					ctr_degree_F_load <= '0';
					ctr_degree_F_rst <= '0';
					reg_degree_G_ce <= '0';
					reg_degree_G_rst <= '0';
					ctr_degree_B_ce <= '0';
					ctr_degree_B_load <= '0';
					ctr_degree_B_rst <= '0';
					sel_ctr_degree_B <= '0';
					reg_degree_C_ce <= '0';
					reg_degree_C_rst <= '0';
					reg_looking_degree_d <= "0";
					reg_looking_degree_ce <= '0';
					reg_swap_ce <= '0';
					reg_swap_rst <= '0';
					sel_address_FB <= '0';
					sel_address_GC <= '0';
					ctr_address_FB_ce <= '1';
					ctr_address_FB_load <= '0';
					ctr_address_GC_ce <= '1';
					ctr_address_GC_load <= '0';
					BC_calculation <= '0';
					enable_external_swap <= '1';
				elsif(degree_F_less_than_degree_G = '1') then
					key_equation_found <= '0';
					signal_inv <= '1';
					sel_new_value_inv <= '1';
					write_enable_FB <= '1';
					write_enable_GC <= '0';
					sel_base_mul <= '0';
					reg_h_ce <= '0';
					ctr_i_ce <= '1';
					ctr_i_load <= '0';
					ctr_i_rst <= '0';
					sel_ctr_i_rst_value <= '0';
					sel_ctr_i_d <= '0';
					reg_j_ce <= '0';
					reg_j_rst <= '0';
					reg_FB_ce <= '0';
					reg_FB_rst <= '0';
					sel_reg_FB <= '0';
					sel_load_new_value_FB <= '0';
					reg_GC_ce <= '0';
					reg_GC_rst <= '0';
					sel_reg_GC <= '0';
					ctr_degree_F_ce <= '0';
					ctr_degree_F_load <= '0';
					ctr_degree_F_rst <= '0';
					reg_degree_G_ce <= '0';
					reg_degree_G_rst <= '0';
					ctr_degree_B_ce <= '0';
					ctr_degree_B_load <= '0';
					ctr_degree_B_rst <= '0';
					sel_ctr_degree_B <= '0';
					reg_degree_C_ce <= '0';
					reg_degree_C_rst <= '0';
					reg_looking_degree_d <= "0";
					reg_looking_degree_ce <= '1';
					reg_swap_ce <= '0';
					reg_swap_rst <= '0';
					sel_address_FB <= '0';
					sel_address_GC <= '0';
					ctr_address_FB_ce <= '1';
					ctr_address_FB_load <= '0';
					ctr_address_GC_ce <= '1';
					ctr_address_GC_load <= '0';
					BC_calculation <= '0';
					enable_external_swap <= '1';
				else
					key_equation_found <= '0';
					signal_inv <= '0';
					sel_new_value_inv <= '0';
					write_enable_FB <= '1';
					write_enable_GC <= '0';
					sel_base_mul <= '0';
					reg_h_ce <= '0';
					ctr_i_ce <= '1';
					ctr_i_load <= '0';
					ctr_i_rst <= '0';
					sel_ctr_i_rst_value <= '0';
					sel_ctr_i_d <= '0';
					reg_j_ce <= '0';
					reg_j_rst <= '0';
					reg_FB_ce <= '0';
					reg_FB_rst <= '0';
					sel_reg_FB <= '0';
					sel_load_new_value_FB <= '0';
					reg_GC_ce <= '0';
					reg_GC_rst <= '0';
					sel_reg_GC <= '0';
					ctr_degree_F_ce <= '0';
					ctr_degree_F_load <= '0';
					ctr_degree_F_rst <= '0';
					reg_degree_G_ce <= '0';
					reg_degree_G_rst <= '0';
					ctr_degree_B_ce <= '0';
					ctr_degree_B_load <= '0';
					ctr_degree_B_rst <= '0';
					sel_ctr_degree_B <= '0';
					reg_degree_C_ce <= '0';
					reg_degree_C_rst <= '0';
					reg_looking_degree_d <= "0";
					reg_looking_degree_ce <= '1';
					reg_swap_ce <= '0';
					reg_swap_rst <= '0';
					sel_address_FB <= '0';
					sel_address_GC <= '0';
					ctr_address_FB_ce <= '1';
					ctr_address_FB_load <= '0';
					ctr_address_GC_ce <= '1';
					ctr_address_GC_load <= '0';
					BC_calculation <= '0';
					enable_external_swap <= '1';
				end if;
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when prepare_i =>
			if(degree_B_equal_degree_C_plus_j = '1') then 
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "1";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			elsif(degree_B_less_than_degree_C_plus_j = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '1';
				ctr_degree_B_load <= '1';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '1';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when finalize_i =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when prepare_load_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when load_B_C =>		
			if(i_minus_j_less_than_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '1';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when mult_add_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '1';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when store_B =>
			if(i_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '0';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '0';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';			
			elsif(reg_looking_degree_q(0) = '1' and FB_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '1';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				sel_new_value_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_load <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= '0';
				sel_ctr_i_d <= '0';
				reg_j_ce <= '0';
				reg_j_rst <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				sel_load_new_value_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				ctr_degree_F_ce <= '0';
				ctr_degree_F_load <= '0';
				ctr_degree_F_rst <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				ctr_degree_B_ce <= '0';
				ctr_degree_B_load <= '0';
				ctr_degree_B_rst <= '0';
				sel_ctr_degree_B <= '0';
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= '0';
				ctr_address_FB_ce <= '1';
				ctr_address_FB_load <= '0';
				ctr_address_GC_ce <= '1';
				ctr_address_GC_load <= '0';
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when prepare_final_swap =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '1';
			ctr_i_load <= '1';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when preparel_swap_address =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when prepare_load_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when load_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when store_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '1';
			ctr_i_load <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '0';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '1';
			ctr_address_FB_load <= '1';
			ctr_address_GC_ce <= '1';
			ctr_address_GC_load <= '1';
			BC_calculation <= '0';
			enable_external_swap <= '0';
		when final =>
			key_equation_found <= '1';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '1';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '1';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '0';
		when others =>
			key_equation_found <= '0';
			signal_inv <= '0';
			sel_new_value_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_load <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= '0';
			sel_ctr_i_d <= '0';
			reg_j_ce <= '0';
			reg_j_rst <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			sel_load_new_value_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			ctr_degree_F_ce <= '0';
			ctr_degree_F_load <= '0';
			ctr_degree_F_rst <= '1';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			ctr_degree_B_ce <= '0';
			ctr_degree_B_load <= '0';
			ctr_degree_B_rst <= '1';
			sel_ctr_degree_B <= '0';
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= '0';
			ctr_address_FB_ce <= '0';
			ctr_address_FB_load <= '0';
			ctr_address_GC_ce <= '0';
			ctr_address_GC_load <= '0';
			BC_calculation <= '0';
			enable_external_swap <= '0';
	end case;
end process;

New_State : process(actual_state, FB_equal_zero, i_equal_zero, i_minus_j_less_than_zero, degree_G_less_equal_final_degree, degree_F_less_than_degree_G,	degree_B_equal_degree_C_plus_j, degree_B_less_than_degree_C_plus_j, reg_looking_degree_q)
begin
	case (actual_state) is
		when reset =>
			next_state <= load_counter;
		when load_counter =>
			next_state <= store_G2t;
		when store_G2t =>
			next_state <= load_first_inv;
		when load_first_inv =>
			next_state <= send_first_inv;
		when send_first_inv =>
			next_state <= prepare_load_F_store_G;
		when prepare_load_F_store_G =>
			next_state <= load_F_store_G;
		when load_F_store_G =>
			next_state <= wait_F;
		when wait_F =>
			if(i_equal_zero = '1') then
				next_state <= prepare_store_B_C;
			else
				next_state <= prepare_load_F_store_G;
			end if;
		when prepare_store_B_C =>
			next_state <= store_B_C;
		when store_B_C =>
			if(i_equal_zero = '1') then
				next_state <= last_store_B_C;
			else
				next_state <= store_B_C;
			end if;
		when last_store_B_C =>
			next_state <= swap_F_G_B_C;
		when swap_F_G_B_C =>
			next_state <= prepare_load_j;
		when prepare_load_j =>
			next_state <= load_j;
		when load_j =>
			next_state <= load_first_G_first_F;
		when load_first_G_first_F =>
			next_state <= load_h;	
		when load_h =>
			next_state <= prepare_load_F_G;
		when prepare_load_F_G =>
			next_state <= load_F_G;
		when load_F_G =>
			next_state <= mult_add_F_G;
		when mult_add_F_G => 
			next_state <= store_F;
		when store_F =>
			if(i_equal_zero = '1') then
				next_state <= prepare_i;
			else
				next_state <= prepare_load_F_G;
			end if;
		when prepare_i =>
			next_state <= finalize_i;
		when finalize_i =>
			next_state <= prepare_load_B_C;
		when prepare_load_B_C =>
			next_state <= load_B_C;
		when load_B_C =>
			next_state <= mult_add_B_C;
		when mult_add_B_C => 	
			next_state <= store_B;
		when store_B =>
			if(i_equal_zero = '1') then
				if(degree_G_less_equal_final_degree = '1') then
					next_state <= prepare_final_swap;
				elsif(degree_F_less_than_degree_G = '1') then
					next_state <= swap_F_G_B_C;
				else
					next_state <= prepare_load_j;
				end if;
			else
				next_state <= prepare_load_B_C;
			end if;
		when prepare_final_swap =>
			next_state <= preparel_swap_address;
		when preparel_swap_address =>
			next_state <= prepare_load_sigma;
		when prepare_load_sigma =>
			next_state <= load_sigma;
		when load_sigma =>
			next_state <= store_sigma;
		when store_sigma =>
			if(i_equal_zero = '1') then
				next_state <= final;
			else
				next_state <= preparel_swap_address;
			end if;
		when final =>
			next_state <= final;
		when others =>
			next_state <= reset;
	end case;
end process;

end Behavioral;

