----------------------------------------------------------------------------------
-- Company: LARC - Escola Politecnica - University of Sao Paulo
-- Engineer: Pedro Maat C. Massolino
-- 
-- Create Date:    05/12/2012 
-- Design Name:    Controller_Solving_Key_Equation_1
-- Module Name:    Controller_Solving_Key_Equation_1
-- Project Name:   McEliece QD-Goppa Decoder
-- Target Devices: Any
-- Tool versions:  Xilinx ISE 13.3 WebPack
--
-- Description: 
-- 
-- The 2nd step in Goppa Code Decoding.
--
-- This is a state machine circuit that controls solving_key_equation_1.
-- This state machine have 3 phases: first phase variable initialization,
-- second computation of polynomial sigma, third step writing the polynomial sigma
-- on a specific memory position.
--
-- This is the first circuit version. It is a non pipeline version of the algorithm, 
-- each coefficient takes more than 1 cycle to be computed.
-- A more optimized version, still non pipeline was made called solving_key_equation_1_v2
-- This improved version, has new address resolution logic and internal degree counters.
--
-- Dependencies: 
--
-- VHDL-93
--
-- Revision: 
-- Revision 1.0
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity controller_solving_key_equation_1 is
	Port (
		clk : in STD_LOGIC;
		rst : in STD_LOGIC;
		ready_inv : in STD_LOGIC;
		FB_equal_zero : in STD_LOGIC;
		i_equal_zero : in STD_LOGIC;
		i_minus_j_less_than_zero : in STD_LOGIC;
		degree_G_less_equal_final_degree : in STD_LOGIC;
		degree_F_less_than_degree_G : in STD_LOGIC;
		degree_B_equal_degree_C_plus_j : in STD_LOGIC;
		degree_B_less_than_degree_C_plus_j : in STD_LOGIC;
		reg_looking_degree_q : in STD_LOGIC_VECTOR(0 downto 0);
		key_equation_found : out STD_LOGIC;
		signal_inv : out STD_LOGIC;
		write_enable_FB : out STD_LOGIC;
		write_enable_GC : out STD_LOGIC;
		sel_base_mul : out STD_LOGIC;
		reg_h_ce : out STD_LOGIC;
		ctr_i_ce : out STD_LOGIC;
		ctr_i_rst : out STD_LOGIC;
		sel_ctr_i_rst_value : out STD_LOGIC_VECTOR(1 downto 0);
		reg_j_ce : out STD_LOGIC;
		reg_FB_ce : out STD_LOGIC;
		reg_FB_rst : out STD_LOGIC;
		sel_reg_FB : out STD_LOGIC;
		reg_GC_ce : out STD_LOGIC;
		reg_GC_rst : out STD_LOGIC;
		sel_reg_GC : out STD_LOGIC;
		reg_degree_F_ce : out STD_LOGIC;
		reg_degree_F_rst : out STD_LOGIC;
		sel_reg_degree_F : out STD_LOGIC;
		reg_degree_G_ce : out STD_LOGIC;
		reg_degree_G_rst : out STD_LOGIC;
		reg_degree_B_ce : out STD_LOGIC;
		reg_degree_B_rst : out STD_LOGIC;
		sel_reg_degree_B : out STD_LOGIC_VECTOR(1 downto 0);
		reg_degree_C_ce : out STD_LOGIC;
		reg_degree_C_rst : out STD_LOGIC;
		reg_looking_degree_d : out STD_LOGIC_VECTOR(0 downto 0);
		reg_looking_degree_ce : out STD_LOGIC;
		reg_swap_ce : out STD_LOGIC;
		reg_swap_rst : out STD_LOGIC;
		sel_int_new_value_FB : out STD_LOGIC;
		sel_address_FB : out STD_LOGIC;
		sel_address_GC : out STD_LOGIC_VECTOR(1 downto 0);
		BC_calculation : out STD_LOGIC;
		enable_external_swap : out STD_LOGIC
	);
end controller_solving_key_equation_1;

architecture Behavioral of controller_solving_key_equation_1 is

type State is (reset, load_counter, store_G2t, prepare_load_F_store_G, load_F_store_G, wait_F, last_load_F_store_G, last_wait_F, store_B_C, last_store_B_C, swap_F_G_B_C, load_j, load_first_G_first_F, send_inv, wait_inv, load_h, prepare_load_F_G, load_F_G, store_F, last_load_F_G, last_store_F, prepare_i, prepare_load_B_C, load_B_C, store_B, last_load_B_C, last_store_B, prepare_final_swap, prepare_load_sigma, load_sigma, last_load_sigma, store_sigma, last_store_sigma, final); 
signal actual_state, next_state : State; 

begin

Clock: process (clk)
begin
	if (clk'event and clk = '1') then
		if (rst = '1') then
			actual_state <= reset;
		else
			actual_state <= next_state;
		end if;        
	end if;
end process;

Output: process(actual_state, ready_inv, FB_equal_zero, i_equal_zero, i_minus_j_less_than_zero, degree_G_less_equal_final_degree, degree_F_less_than_degree_G,	degree_B_equal_degree_C_plus_j, degree_B_less_than_degree_C_plus_j, reg_looking_degree_q)
begin
	case (actual_state) is
		when reset =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '1';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '1';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_counter =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "01";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '1';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '1';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '1';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "01";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when store_G2t =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';			
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "01";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '1';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '1';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "1";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "01";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_F_store_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_F_store_G | last_load_F_store_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when wait_F =>
			if(reg_looking_degree_q(0) = '1' and FB_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '1';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '1';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= "00";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= "00";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when last_wait_F =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';				
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when store_B_C =>
			if(i_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '1';
				sel_base_mul <= '0';
				reg_h_ce <= '0';				
				ctr_i_ce <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '1';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= "00";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '1';
				sel_base_mul <= '0';
				reg_h_ce <= '0';			
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '1';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '0';
				sel_address_FB <= '0';
				sel_address_GC <= "00";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when last_store_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '1';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '1';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when swap_F_G_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '1';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '1';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '1';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '1';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '1';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_j =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "11";
			reg_j_ce <= '1';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '1';
			sel_address_GC <= "01";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_first_G_first_F =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '1';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "01";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when send_inv =>
			key_equation_found <= '0';
			signal_inv <= '1';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when wait_inv =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '1';
			reg_h_ce <= '0';		
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_h =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '1';
			reg_h_ce <= '1';	
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "1";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "10";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_F_G =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= "10";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when load_F_G | last_load_F_G =>
			if(i_minus_j_less_than_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '1';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when store_F =>
			if(reg_looking_degree_q(0) = '1' and FB_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '1';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '1';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '0';
				enable_external_swap <= '1';
			end if;
		when last_store_F =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '1';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '1';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= "10";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_i =>
			if(degree_B_equal_degree_C_plus_j = '1') then 
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '1';
				sel_ctr_i_rst_value <= "10";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "1";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			elsif(degree_B_less_than_degree_C_plus_j = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '1';
				sel_ctr_i_rst_value <= "10";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '1';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "10";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '1';
				sel_ctr_i_rst_value <= "10";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when prepare_load_B_C =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= "10";
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when load_B_C | last_load_B_C =>
			if(i_minus_j_less_than_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '1';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '0';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '0';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '1';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '1';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when store_B =>
			if(reg_looking_degree_q(0) = '1' and FB_equal_zero = '1') then
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '1';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "01";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '0';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			else
				key_equation_found <= '0';
				signal_inv <= '0';
				write_enable_FB <= '1';
				write_enable_GC <= '0';
				sel_base_mul <= '0';
				reg_h_ce <= '0';
				ctr_i_ce <= '1';
				ctr_i_rst <= '0';
				sel_ctr_i_rst_value <= "00";
				reg_j_ce <= '0';
				reg_FB_ce <= '0';
				reg_FB_rst <= '0';
				sel_reg_FB <= '0';
				reg_GC_ce <= '0';
				reg_GC_rst <= '0';
				sel_reg_GC <= '0';
				reg_degree_F_ce <= '0';
				reg_degree_F_rst <= '0';
				sel_reg_degree_F <= '0';
				reg_degree_G_ce <= '0';
				reg_degree_G_rst <= '0';
				reg_degree_B_ce <= '0';
				reg_degree_B_rst <= '0';
				sel_reg_degree_B <= "00";
				reg_degree_C_ce <= '0';
				reg_degree_C_rst <= '0';
				reg_looking_degree_d <= "0";
				reg_looking_degree_ce <= '1';
				reg_swap_ce <= '0';
				reg_swap_rst <= '0';
				sel_int_new_value_FB <= '1';
				sel_address_FB <= '0';
				sel_address_GC <= "10";
				BC_calculation <= '1';
				enable_external_swap <= '1';
			end if;
		when last_store_B =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '1';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '1';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '1';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '1';
			sel_address_FB <= '0';
			sel_address_GC <= "10";
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when prepare_final_swap =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '1';
		when prepare_load_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when load_sigma | last_load_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '1';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '1';
			enable_external_swap <= '1';
		when store_sigma | last_store_sigma =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '1';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '1';
			ctr_i_rst <= '0';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '0';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '0';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '0';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '0';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '0';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '0';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '0';
		when final =>
			key_equation_found <= '1';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '1';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '1';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '1';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '0';
		when others =>
			key_equation_found <= '0';
			signal_inv <= '0';
			write_enable_FB <= '0';
			write_enable_GC <= '0';
			sel_base_mul <= '0';
			reg_h_ce <= '0';
			ctr_i_ce <= '0';
			ctr_i_rst <= '1';
			sel_ctr_i_rst_value <= "00";
			reg_j_ce <= '0';
			reg_FB_ce <= '0';
			reg_FB_rst <= '1';
			sel_reg_FB <= '0';
			reg_GC_ce <= '0';
			reg_GC_rst <= '1';
			sel_reg_GC <= '0';
			reg_degree_F_ce <= '0';
			reg_degree_F_rst <= '1';
			sel_reg_degree_F <= '0';
			reg_degree_G_ce <= '0';
			reg_degree_G_rst <= '1';
			reg_degree_B_ce <= '0';
			reg_degree_B_rst <= '1';
			sel_reg_degree_B <= "00";
			reg_degree_C_ce <= '0';
			reg_degree_C_rst <= '1';
			reg_looking_degree_d <= "0";
			reg_looking_degree_ce <= '0';
			reg_swap_ce <= '0';
			reg_swap_rst <= '0';
			sel_int_new_value_FB <= '0';
			sel_address_FB <= '0';
			sel_address_GC <= "00";
			BC_calculation <= '0';
			enable_external_swap <= '0';
	end case;
end process;

New_State : process(actual_state, ready_inv, FB_equal_zero, i_equal_zero, i_minus_j_less_than_zero, degree_G_less_equal_final_degree, degree_F_less_than_degree_G,	degree_B_equal_degree_C_plus_j, degree_B_less_than_degree_C_plus_j, reg_looking_degree_q)
begin
	case (actual_state) is
		when reset =>
			next_state <= load_counter;
		when load_counter =>
			next_state <= store_G2t;
		when store_G2t =>
			next_state <= prepare_load_F_store_G;
		when prepare_load_F_store_G =>
			if(i_equal_zero = '1') then
				next_state <= last_load_F_store_G;
			else
				next_state <= load_F_store_G;
			end if;
		when load_F_store_G =>
			next_state <= wait_F;
		when wait_F =>
			next_state <= prepare_load_F_store_G;
		when last_load_F_store_G =>
			next_state <= last_wait_F;
		when last_wait_F =>
			next_state <= store_B_C;
		when store_B_C =>
			if(i_equal_zero = '1') then
				next_state <= last_store_B_C;
			else
				next_state <= store_B_C;
			end if;
		when last_store_B_C =>
			next_state <= swap_F_G_B_C;
		when swap_F_G_B_C =>
			next_state <= load_j;
		when load_j =>
			next_state <= load_first_G_first_F;
		when load_first_G_first_F =>
			next_state <= send_inv;	
		when send_inv =>
			next_state <= wait_inv;
		when wait_inv =>
			if(ready_inv = '1') then
				next_state <= load_h;
			else
				next_state <= wait_inv;
			end if;
		when load_h =>
			next_state <= prepare_load_F_G;
		when prepare_load_F_G =>
			if(i_equal_zero = '1') then
				next_state <= last_load_F_G;
			else
				next_state <= load_F_G;
			end if;
		when load_F_G =>
			next_state <= store_F;
		when store_F =>
			next_state <= prepare_load_F_G;
		when last_load_F_G =>
			next_state <= last_store_F;
		when last_store_F =>
			next_state <= prepare_i;
		when prepare_i =>
			next_state <= prepare_load_B_C;
		when prepare_load_B_C =>
			if(i_equal_zero = '1') then
				next_state <= last_load_B_C;
			else
				next_state <= load_B_C;
			end if;
		when load_B_C =>
			next_state <= store_B;
		when store_B =>
			next_state <= prepare_load_B_C;
		when last_load_B_C =>
			next_state <= last_store_B;
		when last_store_B =>
			if(degree_G_less_equal_final_degree = '1') then
				next_state <= prepare_final_swap;
			elsif(degree_F_less_than_degree_G = '1') then
				next_state <= swap_F_G_B_C;
			else
				next_state <= load_j;
			end if;
		when prepare_final_swap =>
			next_state <= prepare_load_sigma;
		when prepare_load_sigma =>
			if(i_equal_zero = '1') then
				next_state <= last_load_sigma;
			else
				next_state <= load_sigma;
			end if;
		when load_sigma =>
			next_state <= store_sigma;
		when last_load_sigma =>
			next_state <= last_store_sigma;
		when store_sigma =>
			next_state <= prepare_load_sigma;
		when last_store_sigma =>
			next_state <= final;
		when final =>
			next_state <= final;
		when others =>
			next_state <= reset;
	end case;
end process;

end Behavioral;

