----------------------------------------------------------------------------------
-- Company: LARC - Escola Politecnica - University of Sao Paulo
-- Engineer: Pedro Maat C. Massolino
-- 
-- Create Date:    05/12/2012 
-- Design Name:    Product_Generator_GF_2_M
-- Module Name:    Product_Generator_GF_2_M
-- Project Name:   GF_2_M Arithmetic
-- Target Devices: Any
-- Tool versions:  Xilinx ISE 13.3 WebPack
--
-- Description: 
--
-- This circuit is part of the GF(2^m) multiplier.
-- This circuit generates the partial product to be latter used in the multiplier.
-- This version is for primitive polynomials present on the software implementation
-- of binary Goppa codes.
--
-- The circuits parameters
--
-- m :
--
-- The size of the field used in this circuit.
--
-- value :
--
-- Used to select the partial product generated by this circuit of
-- o = a * x^(value)
--
-- Dependencies:
-- VHDL-93
--
-- Revision: 
-- Revision 1.0
-- Additional Comments: 
--
----------------------------------------------------------------------------------
architecture Software_POLYNOMIAL of product_generator_gf_2_m is

constant final_value : integer := value mod m;

begin

GF_2_2 : if m = 2 generate -- x^2 + x^1 + 1
	GF_2_2_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_2_P_1 : if final_value = 1 generate
		o <= ( (a(0) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_3 : if m = 3 generate -- x^3 + x^1 + 1
	GF_2_3_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_3_P_1 : if final_value = 1 generate		
		o <= ( a(1) & (a(0) xor a(2)) & a(2) );
	end generate;
	GF_2_3_P_2 : if final_value = 2 generate
		o <= ( (a(0) xor a(2)) & (a(2) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_4 : if m = 4 generate -- x^4 + x^1 + 1
	GF_2_4_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_4_P_1 : if final_value = 1 generate
		o <= ( a(2 downto 1) & (a(0) xor a(3)) & a(3) );
	end generate;
	GF_2_4_P_2 : if final_value = 2 generate
		o <= ( a(1) & (a(0) xor a(3)) & (a(3) xor a(2)) & a(2) );
	end generate;
	GF_2_4_P_3 : if final_value = 3 generate
		o <= ( (a(0) xor a(3)) & (a(3) xor a(2)) & (a(2) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_5 : if m = 5 generate -- x^5 + x^2 + 1
	GF_2_5_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_5_P_1 : if final_value = 1 generate
		o <= ( a(3) & a(2)  & (a(1) xor a(4)) & a(0) & a(4) );
	end generate;
	GF_2_5_P_2 : if final_value = 2 generate
		o <= ( a(2)  & (a(1) xor a(4)) & (a(0) xor a(3)) & a(4) & a(3) );
	end generate;
	GF_2_5_P_3 : if final_value = 3 generate
		o <= ( (a(1) xor a(4)) & (a(0) xor a(3)) & (a(4) xor a(2)) & a(3) & a(2) );
	end generate;
	GF_2_5_P_4 : if final_value = 4 generate
		o <= ( (a(0) xor a(3)) & (a(4) xor a(2)) & (a(3) xor a(1) xor a(4)) & a(2) & (a(1) xor a(4)) );
	end generate;
end generate;

GF_2_6 : if m = 6 generate -- x^6 + x^1 + 1
	GF_2_6_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_6_P_1 : if final_value = 1 generate
		o <= ( a(4) & a(3) & a(2) & a(1) & (a(0) xor a(5)) & a(5) );
	end generate;
	GF_2_6_P_2 : if final_value = 2 generate
		o <= ( a(3) & a(2) & a(1) & (a(0) xor a(5)) & (a(5) xor a(4)) & a(4) );
	end generate;
	GF_2_6_P_3 : if final_value = 3 generate
		o <= ( a(2) & a(1) & (a(0) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & a(3) );
	end generate;
	GF_2_6_P_4 : if final_value = 4 generate
		o <= ( a(1) & (a(0) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & a(2) );
	end generate;
	GF_2_6_P_5 : if final_value = 5 generate
		o <= ( (a(0) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & (a(2) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_7 : if m = 7 generate -- x^7 + x^1 + 1
	GF_2_7_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_7_P_1 : if final_value = 1 generate
		o <= ( a(5) & a(4) & a(3) & a(2) & a(1) & (a(0) xor a(6)) & a(6) );
	end generate;
	GF_2_7_P_2 : if final_value = 2 generate
		o <= ( a(4) & a(3) & a(2) & a(1) & (a(0) xor a(6)) & (a(6) xor a(5)) & a(5) );
	end generate;	
	GF_2_7_P_3 : if final_value = 3 generate
		o <= ( a(3) & a(2) & a(1) & (a(0) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & a(4) );
	end generate;
	GF_2_7_P_4 : if final_value = 4 generate
		o <= ( a(2) & a(1) & (a(0) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & a(3) );
	end generate;
	GF_2_7_P_5 : if final_value = 5 generate
		o <= ( a(1) & (a(0) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & a(2) );
	end generate;
	GF_2_7_P_6 : if final_value = 6 generate
		o <= ( (a(0) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & (a(2) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_8 : if m = 8 generate -- x^8 + x^4 + x^3 + x^2 + 1
	GF_2_8_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_8_P_1 : if final_value = 1 generate
		o <= ( a(6) & a(5) & a(4) & (a(3) xor a(7)) & (a(2) xor a(7)) & (a(1) xor a(7)) & a(0) & a(7) );
	end generate;
	GF_2_8_P_2 : if final_value = 2 generate
		o <= ( a(5) & a(4) & (a(3) xor a(7)) & (a(2) xor a(7) xor a(6)) & (a(1) xor a(7) xor a(6)) & (a(0) xor a(6)) & a(7) & a(6) );
	end generate;
	GF_2_8_P_3 : if final_value = 3 generate
		o <= ( a(4) & (a(3) xor a(7)) & (a(2) xor a(7) xor a(6)) & (a(1) xor a(7) xor a(6) xor a(5)) & (a(0) xor a(6) xor a(5)) & (a(7) xor a(5)) & a(6) & a(5) );
	end generate;
	GF_2_8_P_4 : if final_value = 4 generate
		o <= ( (a(3) xor a(7)) & (a(2) xor a(7) xor a(6)) & (a(1) xor a(7) xor a(6) xor a(5)) & (a(0) xor a(6) xor a(5) xor a(4)) & (a(7) xor a(5) xor a(4)) & (a(6) xor a(4)) & a(5) & a(4) );
	end generate;
	GF_2_8_P_5 : if final_value = 5 generate
		o <= ( (a(2) xor a(7) xor a(6)) & (a(1) xor a(7) xor a(6) xor a(5)) & (a(0) xor a(6) xor a(5) xor a(4)) & (a(5) xor a(4) xor a(3)) & (a(6) xor a(4) xor a(3) xor a(7)) & (a(5) xor a(3) xor a(7)) & a(4) & (a(3) xor a(7)) );
	end generate;
	GF_2_8_P_6 : if final_value = 6 generate
		o <= ( (a(1) xor a(7) xor a(6) xor a(5)) & (a(0) xor a(6) xor a(5) xor a(4)) & (a(5) xor a(4) xor a(3)) & (a(4) xor a(3) xor a(2)) & (a(5) xor a(3) xor a(2) xor a(6)) & (a(4) xor a(2) xor a(7) xor a(6)) & (a(3) xor a(7)) & (a(2) xor a(7) xor a(6)) );
	end generate;
	GF_2_8_P_7 : if final_value = 7 generate
		o <= ( (a(0) xor a(6) xor a(5) xor a(4)) & (a(5) xor a(4) xor a(3)) & (a(4) xor a(3) xor a(2)) & (a(3) xor a(2) xor a(1) xor a(7)) & (a(4) xor a(2) xor a(1) xor a(5)) & (a(3) xor a(1) xor a(6) xor a(5)) & (a(2) xor a(7) xor a(6)) & (a(1) xor a(7) xor a(6) xor a(5)) );
	end generate;
end generate;

GF_2_9 : if m = 9 generate -- x^9 + x^4 + 1
	GF_2_9_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_9_P_1 : if final_value = 1 generate
		o <= ( a(7) & a(6) & a(5) & a(4) & (a(3) xor a(8)) & a(2) & a(1) & a(0) & a(8) );
	end generate;
	GF_2_9_P_2 : if final_value = 2 generate
		o <= ( a(6) & a(5) & a(4) & (a(3) xor a(8)) & (a(2) xor a(7)) & a(1) & a(0) & a(8) & a(7) );
	end generate;
	GF_2_9_P_3 : if final_value = 3 generate
		o <= ( a(5) & a(4) & (a(3) xor a(8)) & (a(2) xor a(7)) & (a(1) xor a(6)) & a(0) & a(8) & a(7) & a(6) );
	end generate;
	GF_2_9_P_4 : if final_value = 4 generate
		o <= ( a(4) & (a(3) xor a(8)) & (a(2) xor a(7)) & (a(1) xor a(6)) & (a(0) xor a(5)) & a(8) & a(7) & a(6) & a(5) );
	end generate;
	GF_2_9_P_5 : if final_value = 5 generate
		o <= ( (a(3) xor a(8)) & (a(2) xor a(7)) & (a(1) xor a(6)) & (a(0) xor a(5)) & (a(8) xor a(4)) & a(7) & a(6) & a(5) & a(4) );
	end generate;
	GF_2_9_P_6 : if final_value = 6 generate
		o <= ( (a(2) xor a(7)) & (a(1) xor a(6)) & (a(0) xor a(5)) & (a(8) xor a(4)) & (a(7) xor a(3) xor a(8)) & a(6) & a(5) & a(4) & (a(3) xor a(8)) );
	end generate;
	GF_2_9_P_7 : if final_value = 7 generate
		o <= ( (a(1) xor a(6)) & (a(0) xor a(5)) & (a(8) xor a(4)) & (a(7) xor a(3) xor a(8)) & (a(6) xor a(2) xor a(7)) & a(5) & a(4) & (a(3) xor a(8)) & (a(2) xor a(7)) );
	end generate;
	GF_2_9_P_8 : if final_value = 8 generate
		o <= ( (a(0) xor a(5)) & (a(8) xor a(4)) & (a(7) xor a(3) xor a(8)) & (a(6) xor a(2) xor a(7)) & (a(5) xor a(1) xor a(6)) & a(4) & (a(3) xor a(8)) & (a(2) xor a(7)) & (a(1) xor a(6)) );
	end generate;
end generate;

GF_2_10 : if m = 10 generate -- x^10 + x^3 + 1
	GF_2_10_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_10_P_1 : if final_value = 1 generate
		o <= ( a(8) & a(7) & a(6) & a(5) & a(4) & a(3) & (a(2) xor a(9)) & a(1) & a(0) & a(9) );
	end generate;
	GF_2_10_P_2 : if final_value = 2 generate
		o <= ( a(7) & a(6) & a(5) & a(4) & a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) & a(0) & a(9) & a(8) );
	end generate;
	GF_2_10_P_3 : if final_value = 3 generate
		o <= ( a(6) & a(5) & a(4) & a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) & (a(0) xor a(7)) & a(9) & a(8) & a(7) );
	end generate;
	GF_2_10_P_4 : if final_value = 4 generate
		o <= ( a(5) & a(4) & a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) & (a(0) xor a(7)) & (a(9) xor a(6)) & a(8) & a(7) & a(6) );
	end generate;
	GF_2_10_P_5 : if final_value = 5 generate
		o <= ( a(4) & a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) & (a(0) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & a(7) & a(6) & a(5) );
	end generate;
	GF_2_10_P_6 : if final_value = 6 generate
		o <= ( a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) & (a(0) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & a(6) & a(5) & a(4) );
	end generate;
	GF_2_10_P_7 : if final_value = 7 generate
		o <= ( (a(2) xor a(9)) & (a(1) xor a(8)) & (a(0) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & a(5) & a(4) & a(3) );
	end generate;
	GF_2_10_P_8 : if final_value = 8 generate
		o <= ( (a(1) xor a(8)) & (a(0) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(9)) & a(4) & a(3) & (a(2) xor a(9)) );
	end generate;
	GF_2_10_P_9 : if final_value = 9 generate
		o <= ( (a(0) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(9)) & (a(4) xor a(1) xor a(8)) & a(3) & (a(2) xor a(9)) & (a(1) xor a(8)) );
	end generate;
end generate;

GF_2_11 : if m = 11 generate -- x^11 + x^2 + 1
	GF_2_11_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_11_P_1 : if final_value = 1 generate
		o <= ( a(9 downto 2) & (a(1) xor a(10)) & a(0) & a(10) );
	end generate;
	GF_2_11_P_2 : if final_value = 2 generate
		o <= ( a(8 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & a(10) & a(9) );
	end generate;
	GF_2_11_P_3 : if final_value = 3 generate
		o <= ( a(7 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & a(9) & a(8) );
	end generate;
	GF_2_11_P_4 : if final_value = 4 generate
		o <= ( a(6 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & a(8) & a(7) );
	end generate;
	GF_2_11_P_5 : if final_value = 5 generate
		o <= ( a(5 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & a(7) & a(6) );
	end generate;
	GF_2_11_P_6 : if final_value = 6 generate
		o <= ( a(4 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & (a(7) xor a(5)) & a(6) & a(5) );
	end generate;
	GF_2_11_P_7 : if final_value = 7 generate
		o <= ( a(3 downto 2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & (a(7) xor a(5)) & (a(6) xor a(4)) & a(5) & a(4) );
	end generate;
	GF_2_11_P_8 : if final_value = 8 generate
		o <= ( a(2) & (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & (a(7) xor a(5)) & (a(6) xor a(4)) & (a(5) xor a(3)) & a(4) & a(3) );
	end generate;
	GF_2_11_P_9 : if final_value = 9 generate
		o <= ( (a(1) xor a(10)) & (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & (a(7) xor a(5)) & (a(6) xor a(4)) & (a(5) xor a(3)) & (a(4) xor a(2)) & a(3) & a(2) );
	end generate;
	GF_2_11_P_10 : if final_value = 10 generate
		o <= ( (a(0) xor a(9)) & (a(10) xor a(8)) & (a(9) xor a(7)) & (a(8) xor a(6)) & (a(7) xor a(5)) & (a(6) xor a(4)) & (a(5) xor a(3)) & (a(4) xor a(2)) & (a(3) xor a(1) xor a(10)) & a(2) & (a(1) xor a(10)) );
	end generate;
end generate;

GF_2_12 : if m = 12 generate -- x^12 + x^6 + x^4 + x^1 + 1
	GF_2_12_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_12_P_1 : if final_value = 1 generate
		o <= ( a(10) & a(9) & a(8) & a(7) & a(6) & (a(5) xor a(11)) & a(4) & (a(3) xor a(11)) & a(2) & a(1) & (a(0) xor a(11)) & a(11) );
	end generate;
	GF_2_12_P_2 : if final_value = 2 generate
		o <= ( a(9) & a(8) & a(7) & a(6) & (a(5) xor a(11)) & (a(4) xor a(10)) & (a(3) xor a(11)) & (a(2) xor a(10)) & a(1) & (a(0) xor a(11)) & (a(11) xor a(10)) & a(10) );
	end generate;
	GF_2_12_P_3 : if final_value = 3 generate
		o <= ( a(8) & a(7) & a(6) & (a(5) xor a(11)) & (a(4) xor a(10)) & (a(3) xor a(11) xor a(9)) & (a(2) xor a(10)) & (a(1) xor a(9)) & (a(0) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & a(9) );
	end generate;
	GF_2_12_P_4 : if final_value = 4 generate
		o <= ( a(7) & a(6) & (a(5) xor a(11)) & (a(4) xor a(10)) & (a(3) xor a(11) xor a(9)) & (a(2) xor a(10) xor a(8)) & (a(1) xor a(9)) & (a(0) xor a(11) xor a(8)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & a(8) );
	end generate;
	GF_2_12_P_5 : if final_value = 5 generate
		o <= ( a(6) & (a(5) xor a(11)) & (a(4) xor a(10)) & (a(3) xor a(11) xor a(9)) & (a(2) xor a(10) xor a(8)) & (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8)) & (a(11) xor a(10) xor a(7)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & a(7) );
	end generate;
	GF_2_12_P_6 : if final_value = 6 generate
		o <= ( (a(5) xor a(11)) & (a(4) xor a(10)) & (a(3) xor a(11) xor a(9)) & (a(2) xor a(10) xor a(8)) & (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8) xor a(6)) & (a(11) xor a(10) xor a(7)) & (a(10) xor a(9) xor a(6)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & a(6) );
	end generate;
	GF_2_12_P_7 : if final_value = 7 generate
		o <= ( (a(4) xor a(10)) & (a(3) xor a(11) xor a(9)) & (a(2) xor a(10) xor a(8)) & (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8) xor a(6)) & (a(10) xor a(7) xor a(5)) & (a(10) xor a(9) xor a(6)) & (a(9) xor a(8) xor a(5) xor a(11)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5) xor a(11)) & (a(5) xor a(11)) );
	end generate;
	GF_2_12_P_8 : if final_value = 8 generate
		o <= ( (a(3) xor a(11) xor a(9)) & (a(2) xor a(10) xor a(8)) & (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8) xor a(6)) & (a(10) xor a(7) xor a(5)) & (a(9) xor a(6) xor a(4)) & (a(9) xor a(8) xor a(5) xor a(11)) & (a(8) xor a(7) xor a(4) xor a(10)) & (a(7) xor a(6)) & (a(6) xor a(5) xor a(11)) & (a(5) xor a(11) xor a(4) xor a(10)) & (a(4) xor a(10)) );
	end generate;
	GF_2_12_P_9 : if final_value = 9 generate
		o <= ( (a(2) xor a(10) xor a(8)) & (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8) xor a(6)) & (a(10) xor a(7) xor a(5)) & (a(9) xor a(6) xor a(4)) & (a(8) xor a(5) xor a(3)) & (a(8) xor a(7) xor a(4) xor a(10)) & (a(7) xor a(6) xor a(3) xor a(11) xor a(9)) & (a(6) xor a(5) xor a(11)) & (a(5) xor a(11) xor a(4) xor a(10)) & (a(4) xor a(10) xor a(3) xor a(11) xor a(9)) & (a(3) xor a(11) xor a(9)) );
	end generate;
	GF_2_12_P_10 : if final_value = 10 generate
		o <= ( (a(1) xor a(9) xor a(7)) & (a(0) xor a(11) xor a(8) xor a(6)) & (a(10) xor a(7) xor a(5)) & (a(9) xor a(6) xor a(4)) & (a(8) xor a(5) xor a(3)) & (a(7) xor a(4) xor a(2)) & (a(7) xor a(6) xor a(3) xor a(11) xor a(9)) & (a(6) xor a(5) xor a(11) xor a(2) xor a(10) xor a(8)) & (a(5) xor a(11) xor a(4) xor a(10)) & (a(4) xor a(10) xor a(3) xor a(11) xor a(9)) & (a(3) xor a(11) xor a(9) xor a(2) xor a(10) xor a(8)) & (a(2) xor a(10) xor a(8)) );
	end generate;
	GF_2_12_P_11 : if final_value = 11 generate
		o <= ( (a(0) xor a(11) xor a(8) xor a(6)) & (a(10) xor a(7) xor a(5)) & (a(9) xor a(6) xor a(4)) & (a(8) xor a(5) xor a(3)) & (a(7) xor a(4) xor a(2)) & (a(6) xor a(3) xor a(11) xor a(1)) & (a(6) xor a(5) xor a(11) xor a(2) xor a(10) xor a(8)) & (a(5) xor a(11) xor a(4) xor a(10) xor a(1) xor a(9) xor a(7)) & (a(4) xor a(10) xor a(3) xor a(11) xor a(9)) & (a(3) xor a(11) xor a(9) xor a(2) xor a(10) xor a(8)) & (a(2) xor a(10) xor a(8) xor a(1) xor a(9) xor a(7)) & (a(1) xor a(9) xor a(7)) );
	end generate;
end generate;

GF_2_13 : if m = 13 generate -- x^13 + x^4 + x^3 + x^1 + 1
	GF_2_13_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_13_P_1 : if final_value = 1 generate
		o <= ( a(11 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12)) & a(1) & (a(0) xor a(12)) & a(12) );
	end generate;
	GF_2_13_P_2 : if final_value = 2 generate
		o <= ( a(10 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11)) & (a(0) xor a(12)) & (a(12) xor a(11)) & a(11) );
	end generate;
	GF_2_13_P_3 : if final_value = 3 generate
		o <= ( a(9 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10)) & (a(12) xor a(11)) & (a(11) xor a(10)) & a(10) );
	end generate;
	GF_2_13_P_4 : if final_value = 4 generate
		o <= ( a(8 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9)) & (a(11) xor a(10)) & (a(10) xor a(9)) & a(9) );
	end generate;
	GF_2_13_P_5 : if final_value = 5 generate
		o <= ( a(7 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8)) & (a(10) xor a(9)) & (a(9) xor a(8)) & a(8) );
	end generate;
	GF_2_13_P_6 : if final_value = 6 generate
		o <= ( a(6 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7)) & (a(9) xor a(8)) & (a(8) xor a(7)) & a(7) );
	end generate;
	GF_2_13_P_7 : if final_value = 7 generate
		o <= ( a(5 downto 4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6)) & (a(8) xor a(7)) & (a(7) xor a(6)) & a(6) );
	end generate;
	GF_2_13_P_8 : if final_value = 8 generate
		o <= ( a(4) & (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6) xor a(5)) & (a(8) xor a(7) xor a(5)) & (a(7) xor a(6)) & (a(6) xor a(5)) & a(5) );
	end generate;
	GF_2_13_P_9 : if final_value = 9 generate
		o <= ( (a(3) xor a(12)) & (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6) xor a(5)) & (a(8) xor a(7) xor a(5) xor a(4)) & (a(7) xor a(6) xor a(4)) & (a(6) xor a(5)) & (a(5) xor a(4)) & a(4) );
	end generate;
	GF_2_13_P_10 : if final_value = 10 generate
		o <= ( (a(2) xor a(12) xor a(11)) & (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6) xor a(5)) & (a(8) xor a(7) xor a(5) xor a(4)) & (a(7) xor a(6) xor a(4) xor a(3) xor a(12)) & (a(6) xor a(5) xor a(3) xor a(12)) & (a(5) xor a(4)) & (a(4) xor a(3) xor a(12)) & (a(3) xor a(12)) );
	end generate;
	GF_2_13_P_11 : if final_value = 11 generate
		o <= ( (a(1) xor a(11) xor a(10)) & (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6) xor a(5)) & (a(8) xor a(7) xor a(5) xor a(4)) & (a(7) xor a(6) xor a(4) xor a(3) xor a(12)) & (a(6) xor a(5) xor a(3) xor a(2) xor a(11)) & (a(5) xor a(4) xor a(2) xor a(12) xor a(11)) & (a(4) xor a(3) xor a(12)) & (a(3) xor a(2) xor a(11)) & (a(2) xor a(12) xor a(11)) );
	end generate;
	GF_2_13_P_12 : if final_value = 12 generate
		o <= ( (a(0) xor a(12) xor a(10) xor a(9)) & (a(12) xor a(11) xor a(9) xor a(8)) & (a(11) xor a(10) xor a(8) xor a(7)) & (a(10) xor a(9) xor a(7) xor a(6)) & (a(9) xor a(8) xor a(6) xor a(5)) & (a(8) xor a(7) xor a(5) xor a(4)) & (a(7) xor a(6) xor a(4) xor a(3) xor a(12)) & (a(6) xor a(5) xor a(3) xor a(2) xor a(11)) & (a(5) xor a(4) xor a(2) xor a(12) xor a(1) xor a(10)) & (a(4) xor a(3) xor a(12) xor a(1) xor a(11) xor a(10)) & (a(3) xor a(2) xor a(11)) & (a(2) xor a(12) xor a(1) xor a(10)) & (a(1) xor a(11) xor a(10)) );
	end generate;
end generate;

GF_2_14 : if m = 14 generate -- x^14 + x^5 + x^3 + x^1 + 1
	GF_2_14_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_14_P_1 : if final_value = 1 generate
		o <= ( a(12) & a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(13)) & a(3) & (a(2) xor a(13)) & a(1) & (a(0) xor a(13)) & a(13) );
	end generate;
	GF_2_14_P_2 : if final_value = 2 generate
		o <= ( a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(13)) & (a(13) xor a(12)) & a(12) );
	end generate;
	GF_2_14_P_3 : if final_value = 3 generate
		o <= ( a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12)) & (a(0) xor a(13) xor a(11)) & (a(13) xor a(12)) & (a(12) xor a(11)) & a(11) );
	end generate;
	GF_2_14_P_4 : if final_value = 4 generate
		o <= ( a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11)) & (a(13) xor a(12) xor a(10)) & (a(12) xor a(11)) & (a(11) xor a(10)) & a(10) );
	end generate;
	GF_2_14_P_5 : if final_value = 5 generate
		o <= ( a(8) & a(7) & a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10)) & (a(12) xor a(11) xor a(9)) & (a(11) xor a(10)) & (a(10) xor a(9)) & a(9) );
	end generate;
	GF_2_14_P_6 : if final_value = 6 generate
		o <= ( a(7) & a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9)) & (a(11) xor a(10) xor a(8)) & (a(10) xor a(9)) & (a(9) xor a(8)) & a(8) );
	end generate;
	GF_2_14_P_7 : if final_value = 7 generate
		o <= ( a(6) & a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8)) & (a(10) xor a(9) xor a(7)) & (a(9) xor a(8)) & (a(8) xor a(7)) & a(7) );
	end generate;
	GF_2_14_P_8 : if final_value = 8 generate
		o <= ( a(5) & (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7)) & (a(9) xor a(8) xor a(6)) & (a(8) xor a(7)) & (a(7) xor a(6)) & a(6) );
	end generate;
	GF_2_14_P_9 : if final_value = 9 generate
		o <= ( (a(4) xor a(13)) & (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7) xor a(5)) & (a(9) xor a(8) xor a(6)) & (a(8) xor a(7) xor a(5)) & (a(7) xor a(6)) & (a(6) xor a(5)) & a(5) );
	end generate;
	GF_2_14_P_10 : if final_value = 10 generate
		o <= ( (a(3) xor a(12)) & (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7) xor a(5)) & (a(9) xor a(8) xor a(6) xor a(4) xor a(13)) & (a(8) xor a(7) xor a(5)) & (a(7) xor a(6) xor a(4) xor a(13)) & (a(6) xor a(5)) & (a(5) xor a(4) xor a(13)) & (a(4) xor a(13)) );
	end generate;
	GF_2_14_P_11 : if final_value = 11 generate
		o <= ( (a(2) xor a(13) xor a(11)) & (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7) xor a(5)) & (a(9) xor a(8) xor a(6) xor a(4) xor a(13)) & (a(8) xor a(7) xor a(5) xor a(3) xor a(12)) & (a(7) xor a(6) xor a(4) xor a(13)) & (a(6) xor a(5) xor a(3) xor a(12)) & (a(5) xor a(4) xor a(13)) & (a(4) xor a(13) xor a(3) xor a(12)) & (a(3) xor a(12)) );
	end generate;
	GF_2_14_P_12 : if final_value = 12 generate
		o <= ( (a(1) xor a(12) xor a(10)) & (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7) xor a(5)) & (a(9) xor a(8) xor a(6) xor a(4) xor a(13)) & (a(8) xor a(7) xor a(5) xor a(3) xor a(12)) & (a(7) xor a(6) xor a(4) xor a(2) xor a(11)) & (a(6) xor a(5) xor a(3) xor a(12)) & (a(5) xor a(4) xor a(2) xor a(11)) & (a(4) xor a(13) xor a(3) xor a(12)) & (a(3) xor a(12) xor a(2) xor a(13) xor a(11)) & (a(2) xor a(13) xor a(11)) );
	end generate;
	GF_2_14_P_13 : if final_value = 13 generate
		o <= ( (a(0) xor a(13) xor a(11) xor a(9)) & (a(13) xor a(12) xor a(10) xor a(8)) & (a(12) xor a(11) xor a(9) xor a(7)) & (a(11) xor a(10) xor a(8) xor a(6)) & (a(10) xor a(9) xor a(7) xor a(5)) & (a(9) xor a(8) xor a(6) xor a(4) xor a(13)) & (a(8) xor a(7) xor a(5) xor a(3) xor a(12)) & (a(7) xor a(6) xor a(4) xor a(2) xor a(11)) & (a(6) xor a(5) xor a(3) xor a(1) xor a(10)) & (a(5) xor a(4) xor a(2) xor a(11)) & (a(4) xor a(13) xor a(3) xor a(1) xor a(10)) & (a(3) xor a(12) xor a(2) xor a(13) xor a(11)) & (a(2) xor a(13) xor a(11) xor a(1) xor a(12) xor a(10)) & (a(1) xor a(12) xor a(10)) );
	end generate;
end generate;

GF_2_15 : if m = 15 generate -- x^15 + x^1 + 1
	GF_2_15_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_15_P_1 : if final_value = 1 generate
		o <= ( a(13 downto 1) & (a(0) xor a(14)) & a(14) );
	end generate;
	GF_2_15_P_2 : if final_value = 2 generate
		o <= ( a(12 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & a(13) );
	end generate;
	GF_2_15_P_3 : if final_value = 3 generate
		o <= ( a(11 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & a(12) );
	end generate;
	GF_2_15_P_4 : if final_value = 4 generate
		o <= ( a(10 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & a(11) );
	end generate;
	GF_2_15_P_5 : if final_value = 5 generate
		o <= ( a(9 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & a(10) );
	end generate;
	GF_2_15_P_6 : if final_value = 6 generate
		o <= ( a(8 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & a(9) );
	end generate;
	GF_2_15_P_7 : if final_value = 7 generate
		o <= ( a(7 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & a(8) );
	end generate;
	GF_2_15_P_8 : if final_value = 8 generate
		o <= ( a(6 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & a(7) );
	end generate;
	GF_2_15_P_9 : if final_value = 9 generate
		o <= ( a(5 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & a(6) );
	end generate;
	GF_2_15_P_10 : if final_value = 10 generate
		o <= ( a(4 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5)) & a(5) );
	end generate;
	GF_2_15_P_11 : if final_value = 11 generate
		o <= ( a(3 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & a(4) );
	end generate;
	GF_2_15_P_12 : if final_value = 12 generate
		o <= ( a(2 downto 1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & a(3) );
	end generate;
	GF_2_15_P_13 : if final_value = 13 generate
		o <= ( a(1) & (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & a(2) );
	end generate;
	GF_2_15_P_14 : if final_value = 14 generate
		o <= ( (a(0) xor a(14)) & (a(14) xor a(13)) & (a(13) xor a(12)) & (a(12) xor a(11)) & (a(11) xor a(10)) & (a(10) xor a(9)) & (a(9) xor a(8)) & (a(8) xor a(7)) & (a(7) xor a(6)) & (a(6) xor a(5)) & (a(5) xor a(4)) & (a(4) xor a(3)) & (a(3) xor a(2)) & (a(2) xor a(1)) & a(1) );
	end generate;
end generate;

GF_2_16 : if m = 16 generate -- x^16 + x^5 + x^3 + x^2 + 1
	GF_2_16_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_16_P_1 : if final_value = 1 generate
		o <= ( a(14) & a(13) & a(12) & a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & a(3) & (a(2) xor a(15)) & (a(1) xor a(15)) & a(0) & a(15) );
	end generate;
	GF_2_16_P_2 : if final_value = 2 generate
		o <= ( a(13) & a(12) & a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15)) & (a(1) xor a(15) xor a(14)) & (a(0) xor a(14)) & a(15) & a(14) );
	end generate;
	GF_2_16_P_3 : if final_value = 3 generate
		o <= ( a(12) & a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14)) & (a(0) xor a(14) xor a(13)) & (a(15) xor a(13)) & a(14) & a(13) );
	end generate;
	GF_2_16_P_4 : if final_value = 4 generate
		o <= ( a(11) & a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13)) & (a(15) xor a(13) xor a(12)) & (a(14) xor a(12)) & a(13) & a(12) );
	end generate;
	GF_2_16_P_5 : if final_value = 5 generate
		o <= ( a(10) & a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12)) & (a(14) xor a(12) xor a(11)) & (a(13) xor a(11)) & a(12) & a(11) );
	end generate;
	GF_2_16_P_6 : if final_value = 6 generate
		o <= ( a(9) & a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11)) & (a(13) xor a(11) xor a(10)) & (a(12) xor a(10)) & a(11) & a(10) );
	end generate;
	GF_2_16_P_7 : if final_value = 7 generate
		o <= ( a(8) & a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10)) & (a(12) xor a(10) xor a(9)) & (a(11) xor a(9)) & a(10) & a(9) );
	end generate;
	GF_2_16_P_8 : if final_value = 8 generate
		o <= ( a(7) & a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9)) & (a(11) xor a(9) xor a(8)) & (a(10) xor a(8)) & a(9) & a(8) );
	end generate;
	GF_2_16_P_9 : if final_value = 9 generate
		o <= ( a(6) & a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8)) & (a(10) xor a(8) xor a(7)) & (a(9) xor a(7)) & a(8) & a(7) );
	end generate;
	GF_2_16_P_10 : if final_value = 10 generate
		o <= ( a(5) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7)) & (a(9) xor a(7) xor a(6)) & (a(8) xor a(6)) & a(7) & a(6) );
	end generate;
	GF_2_16_P_11 : if final_value = 11 generate
		o <= ( (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7) xor a(5)) & (a(9) xor a(7) xor a(6)) & (a(8) xor a(6) xor a(5)) & (a(7) xor a(5)) & a(6) & a(5) );
	end generate;
	GF_2_16_P_12 : if final_value = 12 generate
		o <= ( (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7) xor a(5)) & (a(9) xor a(7) xor a(6) xor a(4) xor a(15)) & (a(8) xor a(6) xor a(5)) & (a(7) xor a(5) xor a(4) xor a(15)) & (a(6) xor a(4) xor a(15)) & a(5) & (a(4) xor a(15)) );
	end generate;
	GF_2_16_P_13 : if final_value = 13 generate
		o <= ( (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7) xor a(5)) & (a(9) xor a(7) xor a(6) xor a(4) xor a(15)) & (a(8) xor a(6) xor a(5) xor a(3) xor a(14)) & (a(7) xor a(5) xor a(4) xor a(15)) & (a(6) xor a(4) xor a(15) xor a(3) xor a(14)) & (a(5) xor a(3) xor a(14)) & (a(4) xor a(15)) & (a(3) xor a(14)) );
	end generate;
	GF_2_16_P_14 : if final_value = 14 generate
		o <= ( (a(1) xor a(15) xor a(14) xor a(12)) & (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7) xor a(5)) & (a(9) xor a(7) xor a(6) xor a(4) xor a(15)) & (a(8) xor a(6) xor a(5) xor a(3) xor a(14)) & (a(7) xor a(5) xor a(4) xor a(2) xor a(13)) & (a(6) xor a(4) xor a(15) xor a(3) xor a(14)) & (a(5) xor a(3) xor a(14) xor a(2) xor a(15) xor a(13)) & (a(4) xor a(2) xor a(13)) & (a(3) xor a(14)) & (a(2) xor a(15) xor a(13)) );
	end generate;
	GF_2_16_P_15 : if final_value = 15 generate
		o <= ( (a(0) xor a(14) xor a(13) xor a(11)) & (a(15) xor a(13) xor a(12) xor a(10)) & (a(14) xor a(12) xor a(11) xor a(9)) & (a(13) xor a(11) xor a(10) xor a(8)) & (a(12) xor a(10) xor a(9) xor a(7)) & (a(11) xor a(9) xor a(8) xor a(6)) & (a(10) xor a(8) xor a(7) xor a(5)) & (a(9) xor a(7) xor a(6) xor a(4) xor a(15)) & (a(8) xor a(6) xor a(5) xor a(3) xor a(14)) & (a(7) xor a(5) xor a(4) xor a(2) xor a(13)) & (a(6) xor a(4) xor a(3) xor a(1) xor a(12)) & (a(5) xor a(3) xor a(14) xor a(2) xor a(15) xor a(13)) & (a(4) xor a(2) xor a(13) xor a(1) xor a(15) xor a(14) xor a(12)) & (a(3) xor a(1) xor a(15) xor a(12)) & (a(2) xor a(15) xor a(13)) & (a(1) xor a(15) xor a(14) xor a(12)) );
	end generate;
end generate;

GF_2_17 : if m = 17 generate -- x^17 + x^3 + 1
	GF_2_17_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_17_P_1 : if final_value = 1 generate
		o <= ( a(15 downto 3) & (a(2) xor a(16)) & a(1) & a(0) & a(16) );
	end generate;
	GF_2_17_P_2 : if final_value = 2 generate
		o <= ( a(14 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & a(0) & a(16) & a(15) );
	end generate;
	GF_2_17_P_3 : if final_value = 3 generate
		o <= ( a(13 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & a(16) & a(15) & a(14) );
	end generate;
	GF_2_17_P_4 : if final_value = 4 generate
		o <= ( a(12 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & a(15) & a(14) & a(13) );
	end generate;
	GF_2_17_P_5 : if final_value = 5 generate
		o <= ( a(11 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & a(14) & a(13) & a(12) );
	end generate;
	GF_2_17_P_6 : if final_value = 6 generate
		o <= ( a(10 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & a(13) & a(12) & a(11) );
	end generate;
	GF_2_17_P_7 : if final_value = 7 generate
		o <= ( a(9 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & a(12) & a(11) & a(10) );
	end generate;
	GF_2_17_P_8 : if final_value = 8 generate
		o <= ( a(8 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & a(11) & a(10) & a(9) );
	end generate;
	GF_2_17_P_9 : if final_value = 9 generate
		o <= ( a(7 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & a(10) & a(9) & a(8) );
	end generate;
	GF_2_17_P_10 : if final_value = 10 generate
		o <= ( a(6 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & a(9) & a(8) & a(7) );
	end generate;
	GF_2_17_P_11 : if final_value = 11 generate
		o <= ( a(5 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & a(8) & a(7) & a(6) );
	end generate;
	GF_2_17_P_12 : if final_value = 12 generate
		o <= ( a(4 downto 3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & a(7) & a(6) & a(5) );
	end generate;
	GF_2_17_P_13 : if final_value = 13 generate
		o <= ( a(3) & (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & a(6) & a(5) & a(4) );
	end generate;
	GF_2_17_P_14 : if final_value = 14 generate
		o <= ( (a(2) xor a(16)) & (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & a(5) & a(4) & a(3) );
	end generate;
	GF_2_17_P_15 : if final_value = 15 generate
		o <= ( (a(1) xor a(15)) & (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(16)) & a(4) & a(3) & (a(2) xor a(16)) );
	end generate;
	GF_2_17_P_16 : if final_value = 16 generate
		o <= ( (a(0) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(16)) & (a(4) xor a(1) xor a(15)) & a(3) & (a(2) xor a(16)) & (a(1) xor a(15)) );
	end generate;
end generate;

GF_2_18 : if m = 18 generate -- x^18 + x^7 + 1
	GF_2_18_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_18_P_1 : if final_value = 1 generate
		o <= ( a(16 downto 7) & (a(6) xor a(17)) & a(5) & a(4) & a(3) & a(2) & a(1) & a(0) & a(17) );
	end generate;
	GF_2_18_P_2 : if final_value = 2 generate
		o <= ( a(15 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & a(4) & a(3) & a(2) & a(1) & a(0) & a(17) & a(16) );
	end generate;
	GF_2_18_P_3 : if final_value = 3 generate
		o <= ( a(14 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & a(3) & a(2) & a(1) & a(0) & a(17) & a(16) & a(15) );
	end generate;
	GF_2_18_P_4 : if final_value = 4 generate
		o <= ( a(13 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & a(2) & a(1) & a(0) & a(17) & a(16) & a(15) & a(14) );
	end generate;
	GF_2_18_P_5 : if final_value = 5 generate
		o <= ( a(12 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & a(1) & a(0) & a(17) & a(16) & a(15) & a(14) & a(13) );
	end generate;
	GF_2_18_P_6 : if final_value = 6 generate
		o <= ( a(11 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & a(0) & a(17) & a(16) & a(15) & a(14) & a(13) & a(12) );
	end generate;
	GF_2_18_P_7 : if final_value = 7 generate
		o <= ( a(10 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & a(17) & a(16) & a(15) & a(14) & a(13) & a(12) & a(11) );
	end generate;
	GF_2_18_P_8 : if final_value = 8 generate
		o <= ( a(9 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & a(16) & a(15) & a(14) & a(13) & a(12) & a(11) & a(10) );
	end generate;
	GF_2_18_P_9 : if final_value = 9 generate
		o <= ( a(8 downto 7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & a(15) & a(14) & a(13) & a(12) & a(11) & a(10) & a(9) );
	end generate;
	GF_2_18_P_10 : if final_value = 10 generate
		o <= ( a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & a(14) & a(13) & a(12) & a(11) & a(10) & a(9) & a(8) );
	end generate;
	GF_2_18_P_11 : if final_value = 11 generate
		o <= ( (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & a(13) & a(12) & a(11) & a(10) & a(9) & a(8) & a(7) );
	end generate;
	GF_2_18_P_12 : if final_value = 12 generate
		o <= ( (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & a(12) & a(11) & a(10) & a(9) & a(8) & a(7) & (a(6) xor a(17)) );
	end generate;
	GF_2_18_P_13 : if final_value = 13 generate
		o <= ( (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & (a(12) xor a(5) xor a(16)) & a(11) & a(10) & a(9) & a(8) & a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) );
	end generate;
	GF_2_18_P_14 : if final_value = 14 generate
		o <= ( (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & (a(12) xor a(5) xor a(16)) & (a(11) xor a(4) xor a(15)) & a(10) & a(9) & a(8) & a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) );
	end generate;
	GF_2_18_P_15 : if final_value = 15 generate
		o <= ( (a(2) xor a(13)) & (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & (a(12) xor a(5) xor a(16)) & (a(11) xor a(4) xor a(15)) & (a(10) xor a(3) xor a(14)) & a(9) & a(8) & a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) );
	end generate;
	GF_2_18_P_16 : if final_value = 16 generate
		o <= ( (a(1) xor a(12)) & (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & (a(12) xor a(5) xor a(16)) & (a(11) xor a(4) xor a(15)) & (a(10) xor a(3) xor a(14)) & (a(9) xor a(2) xor a(13)) & a(8) & a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) );
	end generate;
	GF_2_18_P_17 : if final_value = 17 generate
		o <= ( (a(0) xor a(11)) & (a(17) xor a(10)) & (a(16) xor a(9)) & (a(15) xor a(8)) & (a(14) xor a(7)) & (a(13) xor a(6) xor a(17)) & (a(12) xor a(5) xor a(16)) & (a(11) xor a(4) xor a(15)) & (a(10) xor a(3) xor a(14)) & (a(9) xor a(2) xor a(13)) & (a(8) xor a(1) xor a(12)) & a(7) & (a(6) xor a(17)) & (a(5) xor a(16)) & (a(4) xor a(15)) & (a(3) xor a(14)) & (a(2) xor a(13)) & (a(1) xor a(12)) );
	end generate;
end generate;

GF_2_19 : if m = 19 generate -- x^19 + x^5 + x^2 + x^1 + 1
	GF_2_19_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_19_P_1 : if final_value = 1 generate
		o <= ( a(17 downto 5) & (a(4) xor a(18)) & a(3) & a(2) & (a(1) xor a(18)) & (a(0) xor a(18)) & a(18) );
	end generate;
	GF_2_19_P_2 : if final_value = 2 generate
		o <= ( a(16 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & a(2) & (a(1) xor a(18)) & (a(0) xor a(18) xor a(17)) & (a(18) xor a(17)) & a(17) );
	end generate;
	GF_2_19_P_3 : if final_value = 3 generate
		o <= ( a(15 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18)) & (a(0) xor a(18) xor a(17)) & (a(18) xor a(17) xor a(16)) & (a(17) xor a(16)) & a(16) );
	end generate;
	GF_2_19_P_4 : if final_value = 4 generate
		o <= ( a(14 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17)) & (a(18) xor a(17) xor a(16)) & (a(17) xor a(16) xor a(15)) & (a(16) xor a(15)) & a(15) );
	end generate;
	GF_2_19_P_5 : if final_value = 5 generate
		o <= ( a(13 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16)) & (a(17) xor a(16) xor a(15)) & (a(16) xor a(15) xor a(14)) & (a(15) xor a(14)) & a(14) );
	end generate;
	GF_2_19_P_6 : if final_value = 6 generate
		o <= ( a(12 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15)) & (a(16) xor a(15) xor a(14)) & (a(15) xor a(14) xor a(13)) & (a(14) xor a(13)) & a(13) );
	end generate;
	GF_2_19_P_7 : if final_value = 7 generate
		o <= ( a(11 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14)) & (a(15) xor a(14) xor a(13)) & (a(14) xor a(13) xor a(12)) & (a(13) xor a(12)) & a(12) );
	end generate;
	GF_2_19_P_8 : if final_value = 8 generate
		o <= ( a(10 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13)) & (a(14) xor a(13) xor a(12)) & (a(13) xor a(12) xor a(11)) & (a(12) xor a(11)) & a(11) );
	end generate;
	GF_2_19_P_9 : if final_value = 9 generate
		o <= ( a(9 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12)) & (a(13) xor a(12) xor a(11)) & (a(12) xor a(11) xor a(10)) & (a(11) xor a(10)) & a(10) );
	end generate;
	GF_2_19_P_10 : if final_value = 10 generate
		o <= ( a(8 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11)) & (a(12) xor a(11) xor a(10)) & (a(11) xor a(10) xor a(9)) & (a(10) xor a(9)) & a(9) );
	end generate;
	GF_2_19_P_11 : if final_value = 11 generate
		o <= ( a(7 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10)) & (a(11) xor a(10) xor a(9)) & (a(10) xor a(9) xor a(8)) & (a(9) xor a(8)) & a(8) );
	end generate;
	GF_2_19_P_12 : if final_value = 12 generate
		o <= ( a(6 downto 5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9)) & (a(10) xor a(9) xor a(8)) & (a(9) xor a(8) xor a(7)) & (a(8) xor a(7)) & a(7) );
	end generate;
	GF_2_19_P_13 : if final_value = 13 generate
		o <= ( a(5) & (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8)) & (a(9) xor a(8) xor a(7)) & (a(8) xor a(7) xor a(6)) & (a(7) xor a(6)) & a(6) );
	end generate;
	GF_2_19_P_14 : if final_value = 14 generate
		o <= ( (a(4) xor a(18)) & (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8) xor a(5)) & (a(9) xor a(8) xor a(7)) & (a(8) xor a(7) xor a(6)) & (a(7) xor a(6) xor a(5)) & (a(6) xor a(5)) & a(5) );
	end generate;
	GF_2_19_P_15 : if final_value = 15 generate
		o <= ( (a(3) xor a(17)) & (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8) xor a(5)) & (a(9) xor a(8) xor a(7) xor a(4) xor a(18)) & (a(8) xor a(7) xor a(6)) & (a(7) xor a(6) xor a(5)) & (a(6) xor a(5) xor a(4) xor a(18)) & (a(5) xor a(4) xor a(18)) & (a(4) xor a(18)) );
	end generate;
	GF_2_19_P_16 : if final_value = 16 generate
		o <= ( (a(2) xor a(16)) & (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8) xor a(5)) & (a(9) xor a(8) xor a(7) xor a(4) xor a(18)) & (a(8) xor a(7) xor a(6) xor a(3) xor a(17)) & (a(7) xor a(6) xor a(5)) & (a(6) xor a(5) xor a(4) xor a(18)) & (a(5) xor a(4) xor a(18) xor a(3) xor a(17)) & (a(4) xor a(18) xor a(3) xor a(17)) & (a(3) xor a(17)) );
	end generate;
	GF_2_19_P_17 : if final_value = 17 generate
		o <= ( (a(1) xor a(18) xor a(15)) & (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8) xor a(5)) & (a(9) xor a(8) xor a(7) xor a(4) xor a(18)) & (a(8) xor a(7) xor a(6) xor a(3) xor a(17)) & (a(7) xor a(6) xor a(5) xor a(2) xor a(16)) & (a(6) xor a(5) xor a(4) xor a(18)) & (a(5) xor a(4) xor a(18) xor a(3) xor a(17)) & (a(4) xor a(18) xor a(3) xor a(17) xor a(2) xor a(16)) & (a(3) xor a(17) xor a(2) xor a(16)) & (a(2) xor a(16)) );
	end generate;
	GF_2_19_P_18 : if final_value = 18 generate
		o <= ( (a(0) xor a(18) xor a(17) xor a(14)) & (a(18) xor a(17) xor a(16) xor a(13)) & (a(17) xor a(16) xor a(15) xor a(12)) & (a(16) xor a(15) xor a(14) xor a(11)) & (a(15) xor a(14) xor a(13) xor a(10)) & (a(14) xor a(13) xor a(12) xor a(9)) & (a(13) xor a(12) xor a(11) xor a(8)) & (a(12) xor a(11) xor a(10) xor a(7)) & (a(11) xor a(10) xor a(9) xor a(6)) & (a(10) xor a(9) xor a(8) xor a(5)) & (a(9) xor a(8) xor a(7) xor a(4) xor a(18)) & (a(8) xor a(7) xor a(6) xor a(3) xor a(17)) & (a(7) xor a(6) xor a(5) xor a(2) xor a(16)) & (a(6) xor a(5) xor a(4) xor a(1) xor a(15)) & (a(5) xor a(4) xor a(18) xor a(3) xor a(17)) & (a(4) xor a(18) xor a(3) xor a(17) xor a(2) xor a(16)) & (a(3) xor a(17) xor a(2) xor a(16) xor a(1) xor a(18) xor a(15)) & (a(2) xor a(16) xor a(1) xor a(18) xor a(15)) & (a(1) xor a(18) xor a(15)) );
	end generate;
end generate;

GF_2_20 : if m = 20 generate -- x^20 + x^3 + 1
	GF_2_20_P_0 : if final_value = 0 generate
		o <= a;
	end generate;
	GF_2_20_P_1 : if final_value = 1 generate
		o <= ( a(18 downto 3) & (a(2) xor a(19)) & a(1) & a(0) & a(19) );
	end generate;
	GF_2_20_P_2 : if final_value = 2 generate
		o <= ( a(17 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & a(0) & a(19) & a(18) );
	end generate;
	GF_2_20_P_3 : if final_value = 3 generate
		o <= ( a(16 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & a(19) & a(18) & a(17) );
	end generate;
	GF_2_20_P_4 : if final_value = 4 generate
		o <= ( a(15 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & a(18) & a(17) & a(16) );
	end generate;
	GF_2_20_P_5 : if final_value = 5 generate
		o <= ( a(14 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & a(17) & a(16) & a(15) );
	end generate;
	GF_2_20_P_6 : if final_value = 6 generate
		o <= ( a(13 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & a(16) & a(15) & a(14) );
	end generate;
	GF_2_20_P_7 : if final_value = 7 generate
		o <= ( a(12 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & a(15) & a(14) & a(13) );
	end generate;
	GF_2_20_P_8 : if final_value = 8 generate
		o <= ( a(11 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & a(14) & a(13) & a(12) );
	end generate;
	GF_2_20_P_9 : if final_value = 9 generate
		o <= ( a(10 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & a(13) & a(12) & a(11) );
	end generate;
	GF_2_20_P_10 : if final_value = 10 generate
		o <= ( a(9 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & a(12) & a(11) & a(10) );
	end generate;
	GF_2_20_P_11 : if final_value = 11 generate
		o <= ( a(8 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & a(11) & a(10) & a(9) );
	end generate;
	GF_2_20_P_12 : if final_value = 12 generate
		o <= ( a(7 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & a(10) & a(9) & a(8) );
	end generate;
	GF_2_20_P_13 : if final_value = 13 generate
		o <= ( a(6 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & a(9) & a(8) & a(7) );
	end generate;
	GF_2_20_P_14 : if final_value = 14 generate
		o <= ( a(5 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & a(8) & a(7) & a(6) );
	end generate;
	GF_2_20_P_15 : if final_value = 15 generate
		o <= ( a(4 downto 3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & a(7) & a(6) & a(5) );
	end generate;
	GF_2_20_P_16 : if final_value = 16 generate
		o <= ( a(3) & (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & a(6) & a(5) & a(4) );
	end generate;
	GF_2_20_P_17 : if final_value = 17 generate
		o <= ( (a(2) xor a(19)) & (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & a(5) & a(4) & a(3) );
	end generate;
	GF_2_20_P_18 : if final_value = 18 generate
		o <= ( (a(1) xor a(18)) & (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(19)) & a(4) & a(3) & (a(2) xor a(19)) );
	end generate;
	GF_2_20_P_19 : if final_value = 19 generate
		o <= ( (a(0) xor a(17)) & (a(19) xor a(16)) & (a(18) xor a(15)) & (a(17) xor a(14)) & (a(16) xor a(13)) & (a(15) xor a(12)) & (a(14) xor a(11)) & (a(13) xor a(10)) & (a(12) xor a(9)) & (a(11) xor a(8)) & (a(10) xor a(7)) & (a(9) xor a(6)) & (a(8) xor a(5)) & (a(7) xor a(4)) & (a(6) xor a(3)) & (a(5) xor a(2) xor a(19)) & (a(4) xor a(1) xor a(18)) & a(3) & (a(2) xor a(19)) & (a(1) xor a(18)) );
	end generate;
end generate;

end Software_POLYNOMIAL;

